module andgate(
  input A,       // Input A
  input B,       // Input B
  output Y);     // Output Y
  
  and(Y, A, B);  // Perform logical AND operation on inputs A and B and assign the result to Y
  
endmodule
